// Basic Hello world code
/* 
This code is uses the "$display" to display A basic "Hello World" print to the console.
*/
module hello();
 initial begin
   $display("Hello World");
 end
endmodule
 